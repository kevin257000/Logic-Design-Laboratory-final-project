module board_move(
    input wire [9:0] board_x
);

endmodule